`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/11/03 19:51:55
// Design Name: 
// Module Name: tb_computing_core
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_computing_core();

    //=============================
    // ��������
    //=============================
    parameter WEIGHT_WIDTH = 2048;     // 64*32
    parameter ACT_WIDTH    = 64*448;   // 28672
    parameter RESULT_WIDTH = 8960;     // 64*140 (from design)

    //=============================
    // �ź�����
    //=============================
    reg clk;
    reg [WEIGHT_WIDTH-1:0] i_Weight;
    reg [ACT_WIDTH-1:0]    i_Activation;
    wire [RESULT_WIDTH-1:0] o_result;

    //=============================
    // DUT ʵ����
    //=============================
    computing_core uut (
        .clk(clk),
        .i_Weight(i_Weight),
        .i_Activation(i_Activation),
        .o_result(o_result)
    );

    //=============================
    // ʱ�Ӳ���
    //=============================
    initial begin
        clk = 0;
        forever #5 clk = ~clk; // 100MHz
    end

    //=============================
    // ��������
    //=============================
    integer i;
    reg [31:0] rand_w[0:63];
    reg [447:0] rand_a[0:63];

    // �������������ڴ洢����ʾȨ�ء���������
    reg [31:0] weight_array[0:63];    // 32 bits λ���Ȩ������
    reg [447:0] activation_array[0:63]; // 448 bits λ��ļ�������
    reg [9:0] result_array[0:895];    // 10 bits λ����������

    initial begin
        // ��ʼ��
        i_Weight     = 0;
        i_Activation = 0;

        // ��������ɣ����Զ�Σ�
        for (i = 0; i < 64; i = i + 1) begin
            rand_w[i] = $random;  // 32-bit �����
            rand_a[i] = {$random, $random, $random, $random, $random, $random, $random, $random,
                         $random, $random, $random, $random, $random, $random}; // ƴ��448bit
        end

        // ƴ��Ϊ��������
        for (i = 0; i < 64; i = i + 1) begin
            i_Weight[i*32 +: 32]      = rand_w[i];
            i_Activation[i*448 +: 448] = rand_a[i];
            weight_array[i]           = rand_w[i];               // ���浽Ȩ������
            activation_array[i]       = rand_a[i];               // ���浽��������
        end

        // �Եȼ���ʱ��
        #20;

        // �����ɵڶ���������루��֤��̬�仯��
        for (i = 0; i < 64; i = i + 1) begin
            rand_w[i] = $random;
            rand_a[i] = {$random, $random, $random, $random, $random, $random, $random, $random,
                         $random, $random, $random, $random, $random, $random};
        end

        // ƴ��Ϊ��������
        for (i = 0; i < 64; i = i + 1) begin
            i_Weight[i*32 +: 32]      = rand_w[i];
            i_Activation[i*448 +: 448] = rand_a[i];
            weight_array[i]           = rand_w[i];               // ���浽Ȩ������
            activation_array[i]       = rand_a[i];               // ���浽��������
        end


        #100;
        $finish;
    end

endmodule
