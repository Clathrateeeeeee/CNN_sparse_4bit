`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2025/08/21 10:14:59
// Design Name: 
// Module Name: mult3x3_lut
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


// The function of this code is to multiply the 3b unsigned number by the 3b unsigned number

module mult3x3_lut(
    input       [2:0] a,  // abs(A) lower 3 bits
    input       [2:0] b,  // abs(B) lower 3 bits
    output reg  [5:0] Y
);

    always @(*) 
        begin
            case ({a,b})
                6'b000000: Y = 6'd0;   // 0*0
                6'b000001: Y = 6'd0;   // 0*1
                6'b000010: Y = 6'd0;   // 0*2
                6'b000011: Y = 6'd0;   // 0*3
                6'b000100: Y = 6'd0;   // 0*4
                6'b000101: Y = 6'd0;   // 0*5
                6'b000110: Y = 6'd0;   // 0*6
                6'b000111: Y = 6'd0;   // 0*7

                6'b001000: Y = 6'd0;   // 1*0
                6'b001001: Y = 6'd1;   // 1*1
                6'b001010: Y = 6'd2;   // 1*2
                6'b001011: Y = 6'd3;   // 1*3
                6'b001100: Y = 6'd4;   // 1*4
                6'b001101: Y = 6'd5;   // 1*5
                6'b001110: Y = 6'd6;   // 1*6
                6'b001111: Y = 6'd7;   // 1*7

                6'b010000: Y = 6'd0;   // 2*0
                6'b010001: Y = 6'd2;   // 2*1
                6'b010010: Y = 6'd4;   // 2*2
                6'b010011: Y = 6'd6;   // 2*3
                6'b010100: Y = 6'd8;   // 2*4
                6'b010101: Y = 6'd10;  // 2*5
                6'b010110: Y = 6'd12;  // 2*6
                6'b010111: Y = 6'd14;  // 2*7

                6'b011000: Y = 6'd0;   // 3*0
                6'b011001: Y = 6'd3;   // 3*1
                6'b011010: Y = 6'd6;   // 3*2
                6'b011011: Y = 6'd9;   // 3*3
                6'b011100: Y = 6'd12;  // 3*4
                6'b011101: Y = 6'd15;  // 3*5
                6'b011110: Y = 6'd18;  // 3*6
                6'b011111: Y = 6'd21;  // 3*7

                6'b100000: Y = 6'd0;   // 4*0
                6'b100001: Y = 6'd4;   // 4*1
                6'b100010: Y = 6'd8;   // 4*2
                6'b100011: Y = 6'd12;  // 4*3
                6'b100100: Y = 6'd16;  // 4*4
                6'b100101: Y = 6'd20;  // 4*5
                6'b100110: Y = 6'd24;  // 4*6
                6'b100111: Y = 6'd28;  // 4*7

                6'b101000: Y = 6'd0;   // 5*0
                6'b101001: Y = 6'd5;   // 5*1
                6'b101010: Y = 6'd10;  // 5*2
                6'b101011: Y = 6'd15;  // 5*3
                6'b101100: Y = 6'd20;  // 5*4
                6'b101101: Y = 6'd25;  // 5*5
                6'b101110: Y = 6'd30;  // 5*6
                6'b101111: Y = 6'd35;  // 5*7

                6'b110000: Y = 6'd0;   // 6*0
                6'b110001: Y = 6'd6;   // 6*1
                6'b110010: Y = 6'd12;  // 6*2
                6'b110011: Y = 6'd18;  // 6*3
                6'b110100: Y = 6'd24;  // 6*4
                6'b110101: Y = 6'd30;  // 6*5
                6'b110110: Y = 6'd36;  // 6*6
                6'b110111: Y = 6'd42;  // 6*7

                6'b111000: Y = 6'd0;   // 7*0
                6'b111001: Y = 6'd7;   // 7*1
                6'b111010: Y = 6'd14;  // 7*2
                6'b111011: Y = 6'd21;  // 7*3
                6'b111100: Y = 6'd28;  // 7*4
                6'b111101: Y = 6'd35;  // 7*5
                6'b111110: Y = 6'd42;  // 7*6
                6'b111111: Y = 6'd49;  // 7*7

                default: Y = 6'd0;
            endcase
        end

endmodule


