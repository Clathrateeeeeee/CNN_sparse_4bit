`timescale 1ns/1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/07/17 17:14:38
// Design Name: 
// Module Name: Inbuff
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_ping_pong_ctrl;

    // =================== �������� ===================
    localparam CLK_PERIOD = 10;   // 100 MHz

    // =================== �źŶ��� ===================
    reg  clki;
    reg  rst;
    reg  Ctrl_start;
    reg  done_tile;
    reg  last_tile;
    reg  write_finish;

    wire ping_pong_write;
    wire ping_pong_read;
    wire inbuffer_enout;

    // =================== DUT ���� ===================
    ping_pong_ctrl dut(
        .clki(clki),
        .rst(rst),
        .Ctrl_start(Ctrl_start),
        .done_tile(done_tile),
        .last_tile(last_tile),
        .write_finish(write_finish),
        .ping_pong_write(ping_pong_write),
        .ping_pong_read(ping_pong_read),
        .inbuffer_enout(inbuffer_enout)
    );

    // =================== ʱ�Ӳ��� ===================
    initial begin
        clki = 0;
        forever #(CLK_PERIOD/2) clki = ~clki;
    end

    // =================== ��λ ===================
    initial begin
        rst = 1;
        Ctrl_start = 0;
        done_tile = 0;
        last_tile = 0;
        write_finish = 0;
        #(CLK_PERIOD*5);
        rst = 0;
    end

    // =================== ���񣺲������������� ===================
    task pulse_write_finish;
    begin
        @(posedge clki);
        write_finish <= 1'b1;
        @(posedge clki);
        write_finish <= 1'b0;
    end
    endtask

    task pulse_done_tile;
    begin
        @(posedge clki);
        done_tile <= 1'b1;
        @(posedge clki);
        done_tile <= 1'b0;
    end
    endtask

    // =================== ���� ===================
    initial begin
        // ���� FSM
        #(CLK_PERIOD*10);
        Ctrl_start = 1;
        @(posedge clki);
        Ctrl_start = 0;

        // ---------------- Tile1 ----------------
        // ��д�������
        #(CLK_PERIOD*10);
        pulse_write_finish();

        // ---------------- Tile2 ----------------
        // ģ�� write �� read ��
        #(CLK_PERIOD*20);
        pulse_done_tile();
        #(CLK_PERIOD*10);
        pulse_write_finish();

        // ---------------- Tile3 ----------------
        // ģ�� read �� write ��
        #(CLK_PERIOD*20);
        pulse_write_finish();
        #(CLK_PERIOD*15);
        pulse_done_tile();
        
        #(CLK_PERIOD*20);
        pulse_write_finish();
        #(CLK_PERIOD*15);
        pulse_done_tile();
        
                // ---------------- Tile2 ----------------
        // ģ�� write �� read ��
        #(CLK_PERIOD*20);
        pulse_done_tile();
        #(CLK_PERIOD*10);
        pulse_write_finish();

        // ---------------- Tile3 ----------------
        // ģ�� read �� write ��
        #(CLK_PERIOD*20);
        pulse_write_finish();
        #(CLK_PERIOD*15);
        pulse_done_tile();
        
        #(CLK_PERIOD*20);
        pulse_write_finish();
        #(CLK_PERIOD*15);
        pulse_done_tile();
        
                // ---------------- Tile2 ----------------
        // ģ�� write �� read ��
        #(CLK_PERIOD*20);
        pulse_done_tile();
        #(CLK_PERIOD*10);
        pulse_write_finish();

        // ---------------- Tile3 ----------------
        // ģ�� read �� write ��
        #(CLK_PERIOD*20);
        pulse_write_finish();
        #(CLK_PERIOD*15);
        pulse_done_tile();
        
        #(CLK_PERIOD*20);
        pulse_write_finish();
        #(CLK_PERIOD*15);
        pulse_done_tile();

        // ---------------- ���һ�� tile ----------------
        #(CLK_PERIOD*20);
        last_tile = 1'b1;
        pulse_write_finish();
        #(CLK_PERIOD*20);
        pulse_done_tile();

        #(CLK_PERIOD*50);
        $stop;
    end


endmodule